library verilog;
use verilog.vl_types.all;
entity AluTb is
end AluTb;
